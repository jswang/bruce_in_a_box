module time_averager (
)