-- megafunction wizard: %Shift register (RAM-based)%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTSHIFT_TAPS 

-- ============================================================
-- File Name: ram_shift7.vhd
-- Megafunction Name(s):
-- 			ALTSHIFT_TAPS
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 11.0 Build 157 04/27/2011 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2011 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

ENTITY ram_shift7 IS
	PORT
	(
		clken		: IN STD_LOGIC ;
		clock		: IN STD_LOGIC ;
		shiftin		: IN STD_LOGIC_VECTOR (23 DOWNTO 0);
		shiftout		: OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
		taps		: OUT STD_LOGIC_VECTOR (167 DOWNTO 0)
	);
END ram_shift7;


ARCHITECTURE SYN OF ram_shift7 IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (23 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (167 DOWNTO 0);



	COMPONENT altshift_taps
	GENERIC (
		intended_device_family		: STRING;
		lpm_hint		: STRING;
		lpm_type		: STRING;
		number_of_taps		: NATURAL;
		power_up_state		: STRING;
		tap_distance		: NATURAL;
		width		: NATURAL
	);
	PORT (
			clock	: IN STD_LOGIC ;
			shiftout	: OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
			taps	: OUT STD_LOGIC_VECTOR (167 DOWNTO 0);
			clken	: IN STD_LOGIC ;
			shiftin	: IN STD_LOGIC_VECTOR (23 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	shiftout    <= sub_wire0(23 DOWNTO 0);
	taps    <= sub_wire1(167 DOWNTO 0);

	ALTSHIFT_TAPS_component : ALTSHIFT_TAPS
	GENERIC MAP (
		intended_device_family => "Cyclone IV E",
		lpm_hint => "RAM_BLOCK_TYPE=M4K",
		lpm_type => "altshift_taps",
		number_of_taps => 7,
		power_up_state => "CLEARED",
		tap_distance => 640,
		width => 24
	)
	PORT MAP (
		clock => clock,
		clken => clken,
		shiftin => shiftin,
		shiftout => sub_wire0,
		taps => sub_wire1
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: LPM_HINT STRING "RAM_BLOCK_TYPE=M4K"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altshift_taps"
-- Retrieval info: CONSTANT: NUMBER_OF_TAPS NUMERIC "7"
-- Retrieval info: CONSTANT: POWER_UP_STATE STRING "CLEARED"
-- Retrieval info: CONSTANT: TAP_DISTANCE NUMERIC "640"
-- Retrieval info: CONSTANT: WIDTH NUMERIC "24"
-- Retrieval info: USED_PORT: clken 0 0 0 0 INPUT NODEFVAL "clken"
-- Retrieval info: CONNECT: @clken 0 0 0 0 clken 0 0 0 0
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: USED_PORT: shiftin 0 0 24 0 INPUT NODEFVAL "shiftin[23..0]"
-- Retrieval info: CONNECT: @shiftin 0 0 24 0 shiftin 0 0 24 0
-- Retrieval info: USED_PORT: shiftout 0 0 24 0 OUTPUT NODEFVAL "shiftout[23..0]"
-- Retrieval info: CONNECT: shiftout 0 0 24 0 @shiftout 0 0 24 0
-- Retrieval info: USED_PORT: taps 0 0 168 0 OUTPUT NODEFVAL "taps[167..0]"
-- Retrieval info: CONNECT: taps 0 0 168 0 @taps 0 0 168 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL ram_shift7.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ram_shift7.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ram_shift7.bsf FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ram_shift7_inst.vhd FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ram_shift7.inc FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ram_shift7.cmp FALSE TRUE
-- Retrieval info: LIB_FILE: altera_mf
